--------------------------------------------------------------------------------
--
-- LAB #4
--
--------------------------------------------------------------------------------

Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
Use ieee.std_logic_unsigned.all;

entity ALU is
	Port(	DataIn1: in std_logic_vector(31 downto 0);
		DataIn2: in std_logic_vector(31 downto 0);
		ALUCtrl: in std_logic_vector(4 downto 0);
		Zero: out std_logic;
		ALUResult: out std_logic_vector(31 downto 0) );
end entity ALU;

architecture ALU_Arch of ALU is

	-- ALU components	
	component adder_subtracter
		port(	datain_a: in std_logic_vector(31 downto 0);
			datain_b: in std_logic_vector(31 downto 0);
			add_sub: in std_logic;
			dataout: out std_logic_vector(31 downto 0);
			co: out std_logic);
	end component adder_subtracter;

	component shift_register
		port(	datain: in std_logic_vector(31 downto 0);
		   	dir: in std_logic;
			shamt:	in std_logic_vector(4 downto 0);
			dataout: out std_logic_vector(31 downto 0));
	end component shift_register;

	signal data: std_logic_vector(31 downto 0);
	signal data2: std_logic_vector(31 downto 0);
	signal cout: std_logic_vector(32 downto 0);
	signal co: std_logic;
	signal add_sub: std_logic;

	signal adder: std_logic_vector (31 downto 0);
	signal andi: std_logic_vector(31 downto 0);
	signal ori: std_logic_vector(31 downto 0);
	signal slli: std_logic_vector (31 downto 0);
	signal slri: std_logic_vector (31 downto 0);
	

	

begin
	
	data2 <= DataIn2;
	
	with ALUCtrl(0) select add_sub <=
	'0' when '0',
	'1' when '1',
	'Z' when others; 
	

	A: adder_subtracter port map(DataIn1(31 downto 0), data2(31 downto 0), add_sub, adder(31 downto 0), co);
	andi <= DataIn1 and DataIn2;

	ori <= DataIn1 or DataIn2;
	SL: shift_register port map (DataIn1, '0', DataIn2(4 downto 0), slli); 
	SR: shift_register port map (DataIn1, '1', DataIn2(4 downto 0), slri);

	with ALUCtrl select ALUResult <=
		adder when "00000",
		andi when "00011",
		ori when "00101",
		slli when "00111",
		slri when "01001",
		data2 when "10000",
		"ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ" when others;
		

end architecture ALU_Arch;


